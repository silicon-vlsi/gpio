* Netlist for cascade of three inverters
* MOS model definitions
.model m1 nmos level=3 vto=1v uo=550 vmax=2.0e5
+ cgdo=0.4p cgbo=2.0e-10 cgso=4.0e-11 cjsw=10.e-9
+ mjsw=0.3 tox=1.0e-7 nsub=1.0e16 nfs=1.5e10
+ xj=0.5u ld=0.5u pb=0.75 delta=0.9 eta=0.95
+ kappa=0.45 gamma=0.37

.model p1 pmos level=3 vto=-1v uo=230 vmax=1.9e5
+ cgdo=0.4p cgbo=2.0e-10 cgso=4.0e-11 cjsw=10.e-9
+ mjsw=0.3 tox=1.0e-7 nsub=1.0e16 nfs=1.5e10
+ xj=0.5u ld=0.5u pb=0.75 delta=0.9 eta=0.95
+ kappa=0.45 gamma=0.37
* Subcircuit definition

.subckt inv 1 2 3
m2 2 1 0 0 m1 w=10u l=4u ad=100p pd=40u as=100p
m1 2 1 3 3 p1 w=15u l=4u ad=100p pd=40u as=100p
c1 2 0 0.5p
.ends inv

* Subcircuit calls
x1 1 2 6 inv
x2 2 3 6 inv
x3 3 4 6 inv
cload 4 0 1p

* Electrical source definitions
vdd 6 0 5v
vin 1 0 pulse(0 5 10e-9 5e-9 5e-9 30e-9 50e-9)

* Simulation options & commands
.tran 0.5n 100n uic
.ic v(1)=0
.plot tran v(1) v(2) v(3) v(4)
.print tran v(1) v(2) v(3) v(4)
.option eps=0.5e-3 tnom=50 list node
.end

